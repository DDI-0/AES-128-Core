library ieee;
use ieee.std_logic_1164.all;
use iee.numeric_std.all;

entity aes_fsm is
	po